module bitmap_rom
( input  logic [4:0] char
, input  logic [2:0] row
, input  logic [2:0] col

, output logic       dot
);

    // verilator lint_off ASCRANGE
    logic [0:7] rom [248];
    logic [7:0] addr;

    logic [0:7] data;
    // verilator lint_on ASCRANGE

    assign addr = {char, row};
    assign data = rom[addr];
    assign dot  = data[col];

    initial begin
        // 0
        rom[8'b00000_000] = 8'b00111000;
        rom[8'b00000_001] = 8'b01000100;
        rom[8'b00000_010] = 8'b01001100;
        rom[8'b00000_011] = 8'b01010100;
        rom[8'b00000_100] = 8'b01100100;
        rom[8'b00000_101] = 8'b01000100;
        rom[8'b00000_110] = 8'b00111000;
        rom[8'b00000_111] = 8'b00000000;
        // 1
        rom[8'b00001_000] = 8'b00010000;
        rom[8'b00001_001] = 8'b00110000;
        rom[8'b00001_010] = 8'b01010000;
        rom[8'b00001_011] = 8'b00010000;
        rom[8'b00001_100] = 8'b00010000;
        rom[8'b00001_101] = 8'b00010000;
        rom[8'b00001_110] = 8'b01111100;
        rom[8'b00001_111] = 8'b00000000;
        // 2
        rom[8'b00010_000] = 8'b00111000;
        rom[8'b00010_001] = 8'b01000100;
        rom[8'b00010_010] = 8'b00000100;
        rom[8'b00010_011] = 8'b00001000;
        rom[8'b00010_100] = 8'b00110000;
        rom[8'b00010_101] = 8'b01000000;
        rom[8'b00010_110] = 8'b01111100;
        rom[8'b00010_111] = 8'b00000000;
        // 3
        rom[8'b00011_000] = 8'b00111000;
        rom[8'b00011_001] = 8'b01000100;
        rom[8'b00011_010] = 8'b00000100;
        rom[8'b00011_011] = 8'b00011000;
        rom[8'b00011_100] = 8'b00000100;
        rom[8'b00011_101] = 8'b01000100;
        rom[8'b00011_110] = 8'b00111000;
        rom[8'b00011_111] = 8'b00000000;
        // 4
        rom[8'b00100_000] = 8'b00001000;
        rom[8'b00100_001] = 8'b00011000;
        rom[8'b00100_010] = 8'b00101000;
        rom[8'b00100_011] = 8'b01001000;
        rom[8'b00100_100] = 8'b01111100;
        rom[8'b00100_101] = 8'b00001000;
        rom[8'b00100_110] = 8'b00001000;
        rom[8'b00100_111] = 8'b00000000;
        // 5
        rom[8'b00101_000] = 8'b01111100;
        rom[8'b00101_001] = 8'b01000000;
        rom[8'b00101_010] = 8'b01111000;
        rom[8'b00101_011] = 8'b00000100;
        rom[8'b00101_100] = 8'b00000100;
        rom[8'b00101_101] = 8'b01000100;
        rom[8'b00101_110] = 8'b00111000;
        rom[8'b00101_111] = 8'b00000000;
        // 6
        rom[8'b00110_000] = 8'b00011100;
        rom[8'b00110_001] = 8'b00100000;
        rom[8'b00110_010] = 8'b01000000;
        rom[8'b00110_011] = 8'b01111000;
        rom[8'b00110_100] = 8'b01000100;
        rom[8'b00110_101] = 8'b01000100;
        rom[8'b00110_110] = 8'b00111000;
        rom[8'b00110_111] = 8'b00000000;
        // 7
        rom[8'b00111_000] = 8'b01111100;
        rom[8'b00111_001] = 8'b00000100;
        rom[8'b00111_010] = 8'b00001000;
        rom[8'b00111_011] = 8'b00010000;
        rom[8'b00111_100] = 8'b00100000;
        rom[8'b00111_101] = 8'b00100000;
        rom[8'b00111_110] = 8'b00100000;
        rom[8'b00111_111] = 8'b00000000;
        // 8
        rom[8'b01000_000] = 8'b00111000;
        rom[8'b01000_001] = 8'b01000100;
        rom[8'b01000_010] = 8'b01000100;
        rom[8'b01000_011] = 8'b00111000;
        rom[8'b01000_100] = 8'b01000100;
        rom[8'b01000_101] = 8'b01000100;
        rom[8'b01000_110] = 8'b00111000;
        rom[8'b01000_111] = 8'b00000000;
        // 9
        rom[8'b01001_000] = 8'b00111000;
        rom[8'b01001_001] = 8'b01000100;
        rom[8'b01001_010] = 8'b01000100;
        rom[8'b01001_011] = 8'b00111100;
        rom[8'b01001_100] = 8'b00000100;
        rom[8'b01001_101] = 8'b00001000;
        rom[8'b01001_110] = 8'b01110000;
        rom[8'b01001_111] = 8'b00000000;
        // .
        rom[8'b01010_000] = 8'b00000000;
        rom[8'b01010_001] = 8'b00000000;
        rom[8'b01010_010] = 8'b00000000;
        rom[8'b01010_011] = 8'b00000000;
        rom[8'b01010_100] = 8'b00000000;
        rom[8'b01010_101] = 8'b00000000;
        rom[8'b01010_110] = 8'b00010000;
        rom[8'b01010_111] = 8'b00000000;
        // unk
        rom[8'b01011_000] = 8'b00010001;
        rom[8'b01011_001] = 8'b00100010;
        rom[8'b01011_010] = 8'b01000100;
        rom[8'b01011_011] = 8'b10001000;
        rom[8'b01011_100] = 8'b00010001;
        rom[8'b01011_101] = 8'b00100010;
        rom[8'b01011_110] = 8'b01000100;
        rom[8'b01011_111] = 8'b10001000;
        // P
        rom[8'b01100_000] = 8'b01111100;
        rom[8'b01100_001] = 8'b01000010;
        rom[8'b01100_010] = 8'b01000010;
        rom[8'b01100_011] = 8'b01111100;
        rom[8'b01100_100] = 8'b01000000;
        rom[8'b01100_101] = 8'b01000000;
        rom[8'b01100_110] = 8'b01000000;
        rom[8'b01100_111] = 8'b00000000;
        // r
        rom[8'b01101_000] = 8'b00000000;
        rom[8'b01101_001] = 8'b00000000;
        rom[8'b01101_010] = 8'b01011100;
        rom[8'b01101_011] = 8'b01100000;
        rom[8'b01101_100] = 8'b01000000;
        rom[8'b01101_101] = 8'b01000000;
        rom[8'b01101_110] = 8'b01000000;
        rom[8'b01101_111] = 8'b00000000;
        // e
        rom[8'b01110_000] = 8'b00000000;
        rom[8'b01110_001] = 8'b00000000;
        rom[8'b01110_010] = 8'b00111000;
        rom[8'b01110_011] = 8'b01000100;
        rom[8'b01110_100] = 8'b01111100;
        rom[8'b01110_101] = 8'b01000000;
        rom[8'b01110_110] = 8'b00111000;
        rom[8'b01110_111] = 8'b00000000;
        // s
        rom[8'b01111_000] = 8'b00000000;
        rom[8'b01111_001] = 8'b00000000;
        rom[8'b01111_010] = 8'b00111100;
        rom[8'b01111_011] = 8'b01000000;
        rom[8'b01111_100] = 8'b00111000;
        rom[8'b01111_101] = 8'b00000100;
        rom[8'b01111_110] = 8'b01111000;
        rom[8'b01111_111] = 8'b00000000;
        // b
        rom[8'b10000_000] = 8'b01000000;
        rom[8'b10000_001] = 8'b01000000;
        rom[8'b10000_010] = 8'b01111000;
        rom[8'b10000_011] = 8'b01000100;
        rom[8'b10000_100] = 8'b01000100;
        rom[8'b10000_101] = 8'b01000100;
        rom[8'b10000_110] = 8'b01111000;
        rom[8'b10000_111] = 8'b00000000;
        // u
        rom[8'b10001_000] = 8'b00000000;
        rom[8'b10001_001] = 8'b00000000;
        rom[8'b10001_010] = 8'b01000100;
        rom[8'b10001_011] = 8'b01000100;
        rom[8'b10001_100] = 8'b01000100;
        rom[8'b10001_101] = 8'b01000100;
        rom[8'b10001_110] = 8'b00111000;
        rom[8'b10001_111] = 8'b00000000;
        // t
        rom[8'b10010_000] = 8'b00100000;
        rom[8'b10010_001] = 8'b00100000;
        rom[8'b10010_010] = 8'b01111000;
        rom[8'b10010_011] = 8'b00100000;
        rom[8'b10010_100] = 8'b00100000;
        rom[8'b10010_101] = 8'b00100100;
        rom[8'b10010_110] = 8'b00011000;
        rom[8'b10010_111] = 8'b00000000;
        // o
        rom[8'b10011_000] = 8'b00000000;
        rom[8'b10011_001] = 8'b00000000;
        rom[8'b10011_010] = 8'b00111000;
        rom[8'b10011_011] = 8'b01000100;
        rom[8'b10011_100] = 8'b01000100;
        rom[8'b10011_101] = 8'b01000100;
        rom[8'b10011_110] = 8'b00111000;
        rom[8'b10011_111] = 8'b00000000;
        // n
        rom[8'b10100_000] = 8'b00000000;
        rom[8'b10100_001] = 8'b00000000;
        rom[8'b10100_010] = 8'b01111000;
        rom[8'b10100_011] = 8'b01000100;
        rom[8'b10100_100] = 8'b01000100;
        rom[8'b10100_101] = 8'b01000100;
        rom[8'b10100_110] = 8'b01000100;
        rom[8'b10100_111] = 8'b00000000;
        // a
        rom[8'b10101_000] = 8'b00000000;
        rom[8'b10101_001] = 8'b00000000;
        rom[8'b10101_010] = 8'b00111000;
        rom[8'b10101_011] = 8'b00000100;
        rom[8'b10101_100] = 8'b00111100;
        rom[8'b10101_101] = 8'b01000100;
        rom[8'b10101_110] = 8'b00111100;
        rom[8'b10101_111] = 8'b00000000;
        // W
        rom[8'b10110_000] = 8'b01000010;
        rom[8'b10110_001] = 8'b01000010;
        rom[8'b10110_010] = 8'b01000010;
        rom[8'b10110_011] = 8'b01000010;
        rom[8'b10110_100] = 8'b01011010;
        rom[8'b10110_101] = 8'b01100110;
        rom[8'b10110_110] = 8'b01000010;
        rom[8'b10110_111] = 8'b00000000;
        // i
        rom[8'b10111_000] = 8'b00010000;
        rom[8'b10111_001] = 8'b00000000;
        rom[8'b10111_010] = 8'b00110000;
        rom[8'b10111_011] = 8'b00010000;
        rom[8'b10111_100] = 8'b00010000;
        rom[8'b10111_101] = 8'b00010000;
        rom[8'b10111_110] = 8'b00111000;
        rom[8'b10111_111] = 8'b00000000;
        // M
        rom[8'b11000_000] = 8'b01000010;
        rom[8'b11000_001] = 8'b01100110;
        rom[8'b11000_010] = 8'b01011010;
        rom[8'b11000_011] = 8'b01000010;
        rom[8'b11000_100] = 8'b01000010;
        rom[8'b11000_101] = 8'b01000010;
        rom[8'b11000_110] = 8'b01000010;
        rom[8'b11000_111] = 8'b00000000;
        // L
        rom[8'b11001_000] = 8'b01000000;
        rom[8'b11001_001] = 8'b01000000;
        rom[8'b11001_010] = 8'b01000000;
        rom[8'b11001_011] = 8'b01000000;
        rom[8'b11001_100] = 8'b01000000;
        rom[8'b11001_101] = 8'b01000000;
        rom[8'b11001_110] = 8'b01111110;
        rom[8'b11001_111] = 8'b00000000;
        // :
        rom[8'b11010_000] = 8'b00000000;
        rom[8'b11010_001] = 8'b00000000;
        rom[8'b11010_010] = 8'b00010000;
        rom[8'b11010_011] = 8'b00000000;
        rom[8'b11010_100] = 8'b00000000;
        rom[8'b11010_101] = 8'b00010000;
        rom[8'b11010_110] = 8'b00000000;
        rom[8'b11010_111] = 8'b00000000;
        // B
        rom[8'b11011_000] = 8'b01111100;
        rom[8'b11011_001] = 8'b01000010;
        rom[8'b11011_010] = 8'b01000010;
        rom[8'b11011_011] = 8'b01111100;
        rom[8'b11011_100] = 8'b01000010;
        rom[8'b11011_101] = 8'b01000010;
        rom[8'b11011_110] = 8'b01111100;
        rom[8'b11011_111] = 8'b00000000;
        // micro
        rom[8'b11100_000] = 8'b00000000;
        rom[8'b11100_001] = 8'b00000000;
        rom[8'b11100_010] = 8'b00100010;
        rom[8'b11100_011] = 8'b00100010;
        rom[8'b11100_100] = 8'b00100010;
        rom[8'b11100_101] = 8'b00111100;
        rom[8'b11100_110] = 8'b00100000;
        rom[8'b11100_111] = 8'b01000000;
        // m
        rom[8'b11101_000] = 8'b00000000;
        rom[8'b11101_001] = 8'b00000000;
        rom[8'b11101_010] = 8'b01101000;
        rom[8'b11101_011] = 8'b01010100;
        rom[8'b11101_100] = 8'b01010100;
        rom[8'b11101_101] = 8'b01010100;
        rom[8'b11101_110] = 8'b01010100;
        rom[8'b11101_111] = 8'b00000000;
        // H
        rom[8'b11110_000] = 8'b01000010;
        rom[8'b11110_001] = 8'b01000010;
        rom[8'b11110_010] = 8'b01000010;
        rom[8'b11110_011] = 8'b01111110;
        rom[8'b11110_100] = 8'b01000010;
        rom[8'b11110_101] = 8'b01000010;
        rom[8'b11110_110] = 8'b01000010;
        rom[8'b11110_111] = 8'b00000000;
    end

endmodule : bitmap_rom
