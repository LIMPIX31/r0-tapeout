module bitmap_rom #
( parameter int unsigned ADDR_WIDTH = 6
)
( input  logic [ADDR_WIDTH-1:0] char
, input  logic [2:0] row
, input  logic [2:0] col

, output logic       dot
);

    logic [7:0] rom [1 << (ADDR_WIDTH + 3)];

    logic [ADDR_WIDTH+2:0] addr;

    logic [7:0] data;

    assign addr = {char, row};
    assign data = rom[addr];
    assign dot  = data[col];

    initial begin
        (* font_start *);

        // '.' => 6'b001010
        // ':' => 6'b001011
        // 'B' => 6'b001100
        // 'H' => 6'b001101
        // 'L' => 6'b001110
        // 'M' => 6'b001111
        // 'P' => 6'b010000
        // 'R' => 6'b010001
        // 'a' => 6'b010010
        // 'b' => 6'b010011
        // 'd' => 6'b010100
        // 'e' => 6'b010101
        // 'i' => 6'b010110
        // 'm' => 6'b010111
        // 'n' => 6'b011000
        // 'o' => 6'b011001
        // 'r' => 6'b011010
        // 's' => 6'b011011
        // 't' => 6'b011100
        // 'u' => 6'b011101
        // 'y' => 6'b011110
        // '»' => 6'b011111
        // 'ö' => 6'b100000

        rom[9'b000000_111] = 8'b00000000;
        rom[9'b000000_110] = 8'b00011100;
        rom[9'b000000_101] = 8'b00100010;
        rom[9'b000000_100] = 8'b00100110;
        rom[9'b000000_011] = 8'b00101010;
        rom[9'b000000_010] = 8'b00110010;
        rom[9'b000000_001] = 8'b00100010;
        rom[9'b000000_000] = 8'b00011100;

        rom[9'b000001_111] = 8'b00000000;
        rom[9'b000001_110] = 8'b00111110;
        rom[9'b000001_101] = 8'b00001000;
        rom[9'b000001_100] = 8'b00001000;
        rom[9'b000001_011] = 8'b00001000;
        rom[9'b000001_010] = 8'b00001010;
        rom[9'b000001_001] = 8'b00001100;
        rom[9'b000001_000] = 8'b00001000;

        rom[9'b000010_111] = 8'b00000000;
        rom[9'b000010_110] = 8'b00111110;
        rom[9'b000010_101] = 8'b00000010;
        rom[9'b000010_100] = 8'b00001100;
        rom[9'b000010_011] = 8'b00010000;
        rom[9'b000010_010] = 8'b00100000;
        rom[9'b000010_001] = 8'b00100010;
        rom[9'b000010_000] = 8'b00011100;

        rom[9'b000011_111] = 8'b00000000;
        rom[9'b000011_110] = 8'b00011100;
        rom[9'b000011_101] = 8'b00100010;
        rom[9'b000011_100] = 8'b00100000;
        rom[9'b000011_011] = 8'b00011000;
        rom[9'b000011_010] = 8'b00100000;
        rom[9'b000011_001] = 8'b00100010;
        rom[9'b000011_000] = 8'b00011100;

        rom[9'b000100_111] = 8'b00000000;
        rom[9'b000100_110] = 8'b00010000;
        rom[9'b000100_101] = 8'b00010000;
        rom[9'b000100_100] = 8'b00111110;
        rom[9'b000100_011] = 8'b00010010;
        rom[9'b000100_010] = 8'b00010100;
        rom[9'b000100_001] = 8'b00011000;
        rom[9'b000100_000] = 8'b00010000;

        rom[9'b000101_111] = 8'b00000000;
        rom[9'b000101_110] = 8'b00011100;
        rom[9'b000101_101] = 8'b00100010;
        rom[9'b000101_100] = 8'b00100000;
        rom[9'b000101_011] = 8'b00100000;
        rom[9'b000101_010] = 8'b00011110;
        rom[9'b000101_001] = 8'b00000010;
        rom[9'b000101_000] = 8'b00111110;

        rom[9'b000110_111] = 8'b00000000;
        rom[9'b000110_110] = 8'b00011100;
        rom[9'b000110_101] = 8'b00100010;
        rom[9'b000110_100] = 8'b00100010;
        rom[9'b000110_011] = 8'b00011110;
        rom[9'b000110_010] = 8'b00000010;
        rom[9'b000110_001] = 8'b00000100;
        rom[9'b000110_000] = 8'b00111000;

        rom[9'b000111_111] = 8'b00000000;
        rom[9'b000111_110] = 8'b00000100;
        rom[9'b000111_101] = 8'b00000100;
        rom[9'b000111_100] = 8'b00000100;
        rom[9'b000111_011] = 8'b00001000;
        rom[9'b000111_010] = 8'b00010000;
        rom[9'b000111_001] = 8'b00100000;
        rom[9'b000111_000] = 8'b00111110;

        rom[9'b001000_111] = 8'b00000000;
        rom[9'b001000_110] = 8'b00011100;
        rom[9'b001000_101] = 8'b00100010;
        rom[9'b001000_100] = 8'b00100010;
        rom[9'b001000_011] = 8'b00011100;
        rom[9'b001000_010] = 8'b00100010;
        rom[9'b001000_001] = 8'b00100010;
        rom[9'b001000_000] = 8'b00011100;

        rom[9'b001001_111] = 8'b00000000;
        rom[9'b001001_110] = 8'b00001110;
        rom[9'b001001_101] = 8'b00010000;
        rom[9'b001001_100] = 8'b00100000;
        rom[9'b001001_011] = 8'b00111100;
        rom[9'b001001_010] = 8'b00100010;
        rom[9'b001001_001] = 8'b00100010;
        rom[9'b001001_000] = 8'b00011100;

        rom[9'b001010_111] = 8'b00000000;
        rom[9'b001010_110] = 8'b00001000;
        rom[9'b001010_101] = 8'b00000000;
        rom[9'b001010_100] = 8'b00000000;
        rom[9'b001010_011] = 8'b00000000;
        rom[9'b001010_010] = 8'b00000000;
        rom[9'b001010_001] = 8'b00000000;
        rom[9'b001010_000] = 8'b00000000;

        rom[9'b001011_111] = 8'b00000000;
        rom[9'b001011_110] = 8'b00000000;
        rom[9'b001011_101] = 8'b00001000;
        rom[9'b001011_100] = 8'b00000000;
        rom[9'b001011_011] = 8'b00000000;
        rom[9'b001011_010] = 8'b00001000;
        rom[9'b001011_001] = 8'b00000000;
        rom[9'b001011_000] = 8'b00000000;

        rom[9'b001100_111] = 8'b00000000;
        rom[9'b001100_110] = 8'b00111110;
        rom[9'b001100_101] = 8'b01000010;
        rom[9'b001100_100] = 8'b01000010;
        rom[9'b001100_011] = 8'b00111110;
        rom[9'b001100_010] = 8'b01000010;
        rom[9'b001100_001] = 8'b01000010;
        rom[9'b001100_000] = 8'b00111110;

        rom[9'b001101_111] = 8'b00000000;
        rom[9'b001101_110] = 8'b01000010;
        rom[9'b001101_101] = 8'b01000010;
        rom[9'b001101_100] = 8'b01000010;
        rom[9'b001101_011] = 8'b01111110;
        rom[9'b001101_010] = 8'b01000010;
        rom[9'b001101_001] = 8'b01000010;
        rom[9'b001101_000] = 8'b01000010;

        rom[9'b001110_111] = 8'b00000000;
        rom[9'b001110_110] = 8'b01111110;
        rom[9'b001110_101] = 8'b00000010;
        rom[9'b001110_100] = 8'b00000010;
        rom[9'b001110_011] = 8'b00000010;
        rom[9'b001110_010] = 8'b00000010;
        rom[9'b001110_001] = 8'b00000010;
        rom[9'b001110_000] = 8'b00000010;

        rom[9'b001111_111] = 8'b00000000;
        rom[9'b001111_110] = 8'b01000010;
        rom[9'b001111_101] = 8'b01000010;
        rom[9'b001111_100] = 8'b01000010;
        rom[9'b001111_011] = 8'b01000010;
        rom[9'b001111_010] = 8'b01011010;
        rom[9'b001111_001] = 8'b01100110;
        rom[9'b001111_000] = 8'b01000010;

        rom[9'b010000_111] = 8'b00000000;
        rom[9'b010000_110] = 8'b00000010;
        rom[9'b010000_101] = 8'b00000010;
        rom[9'b010000_100] = 8'b00000010;
        rom[9'b010000_011] = 8'b00111110;
        rom[9'b010000_010] = 8'b01000010;
        rom[9'b010000_001] = 8'b01000010;
        rom[9'b010000_000] = 8'b00111110;

        rom[9'b010001_111] = 8'b00000000;
        rom[9'b010001_110] = 8'b01000010;
        rom[9'b010001_101] = 8'b00100010;
        rom[9'b010001_100] = 8'b00010010;
        rom[9'b010001_011] = 8'b00111110;
        rom[9'b010001_010] = 8'b01000010;
        rom[9'b010001_001] = 8'b01000010;
        rom[9'b010001_000] = 8'b00111110;

        rom[9'b010010_111] = 8'b00000000;
        rom[9'b010010_110] = 8'b00111100;
        rom[9'b010010_101] = 8'b00100010;
        rom[9'b010010_100] = 8'b00111100;
        rom[9'b010010_011] = 8'b00100000;
        rom[9'b010010_010] = 8'b00011100;
        rom[9'b010010_001] = 8'b00000000;
        rom[9'b010010_000] = 8'b00000000;

        rom[9'b010011_111] = 8'b00000000;
        rom[9'b010011_110] = 8'b00011110;
        rom[9'b010011_101] = 8'b00100010;
        rom[9'b010011_100] = 8'b00100010;
        rom[9'b010011_011] = 8'b00100010;
        rom[9'b010011_010] = 8'b00011110;
        rom[9'b010011_001] = 8'b00000010;
        rom[9'b010011_000] = 8'b00000010;

        rom[9'b010100_111] = 8'b00000000;
        rom[9'b010100_110] = 8'b00111100;
        rom[9'b010100_101] = 8'b00100010;
        rom[9'b010100_100] = 8'b00100010;
        rom[9'b010100_011] = 8'b00100010;
        rom[9'b010100_010] = 8'b00111100;
        rom[9'b010100_001] = 8'b00100000;
        rom[9'b010100_000] = 8'b00100000;

        rom[9'b010101_111] = 8'b00000000;
        rom[9'b010101_110] = 8'b00011100;
        rom[9'b010101_101] = 8'b00000010;
        rom[9'b010101_100] = 8'b00111110;
        rom[9'b010101_011] = 8'b00100010;
        rom[9'b010101_010] = 8'b00011100;
        rom[9'b010101_001] = 8'b00000000;
        rom[9'b010101_000] = 8'b00000000;

        rom[9'b010110_111] = 8'b00000000;
        rom[9'b010110_110] = 8'b00011100;
        rom[9'b010110_101] = 8'b00001000;
        rom[9'b010110_100] = 8'b00001000;
        rom[9'b010110_011] = 8'b00001000;
        rom[9'b010110_010] = 8'b00001100;
        rom[9'b010110_001] = 8'b00000000;
        rom[9'b010110_000] = 8'b00001000;

        rom[9'b010111_111] = 8'b00000000;
        rom[9'b010111_110] = 8'b00101010;
        rom[9'b010111_101] = 8'b00101010;
        rom[9'b010111_100] = 8'b00101010;
        rom[9'b010111_011] = 8'b00101010;
        rom[9'b010111_010] = 8'b00010110;
        rom[9'b010111_001] = 8'b00000000;
        rom[9'b010111_000] = 8'b00000000;

        rom[9'b011000_111] = 8'b00000000;
        rom[9'b011000_110] = 8'b00100010;
        rom[9'b011000_101] = 8'b00100010;
        rom[9'b011000_100] = 8'b00100010;
        rom[9'b011000_011] = 8'b00100010;
        rom[9'b011000_010] = 8'b00011110;
        rom[9'b011000_001] = 8'b00000000;
        rom[9'b011000_000] = 8'b00000000;

        rom[9'b011001_111] = 8'b00000000;
        rom[9'b011001_110] = 8'b00011100;
        rom[9'b011001_101] = 8'b00100010;
        rom[9'b011001_100] = 8'b00100010;
        rom[9'b011001_011] = 8'b00100010;
        rom[9'b011001_010] = 8'b00011100;
        rom[9'b011001_001] = 8'b00000000;
        rom[9'b011001_000] = 8'b00000000;

        rom[9'b011010_111] = 8'b00000000;
        rom[9'b011010_110] = 8'b00000010;
        rom[9'b011010_101] = 8'b00000010;
        rom[9'b011010_100] = 8'b00000010;
        rom[9'b011010_011] = 8'b00000110;
        rom[9'b011010_010] = 8'b00111010;
        rom[9'b011010_001] = 8'b00000000;
        rom[9'b011010_000] = 8'b00000000;

        rom[9'b011011_111] = 8'b00000000;
        rom[9'b011011_110] = 8'b00011110;
        rom[9'b011011_101] = 8'b00100000;
        rom[9'b011011_100] = 8'b00011100;
        rom[9'b011011_011] = 8'b00000010;
        rom[9'b011011_010] = 8'b00111100;
        rom[9'b011011_001] = 8'b00000000;
        rom[9'b011011_000] = 8'b00000000;

        rom[9'b011100_111] = 8'b00000000;
        rom[9'b011100_110] = 8'b00011000;
        rom[9'b011100_101] = 8'b00100100;
        rom[9'b011100_100] = 8'b00000100;
        rom[9'b011100_011] = 8'b00000100;
        rom[9'b011100_010] = 8'b00011110;
        rom[9'b011100_001] = 8'b00000100;
        rom[9'b011100_000] = 8'b00000100;

        rom[9'b011101_111] = 8'b00000000;
        rom[9'b011101_110] = 8'b00011100;
        rom[9'b011101_101] = 8'b00100010;
        rom[9'b011101_100] = 8'b00100010;
        rom[9'b011101_011] = 8'b00100010;
        rom[9'b011101_010] = 8'b00100010;
        rom[9'b011101_001] = 8'b00000000;
        rom[9'b011101_000] = 8'b00000000;

        rom[9'b011110_111] = 8'b00011100;
        rom[9'b011110_110] = 8'b00100000;
        rom[9'b011110_101] = 8'b00111100;
        rom[9'b011110_100] = 8'b00100010;
        rom[9'b011110_011] = 8'b00100010;
        rom[9'b011110_010] = 8'b00100010;
        rom[9'b011110_001] = 8'b00000000;
        rom[9'b011110_000] = 8'b00000000;

        rom[9'b011111_111] = 8'b00000010;
        rom[9'b011111_110] = 8'b00000100;
        rom[9'b011111_101] = 8'b00111100;
        rom[9'b011111_100] = 8'b01000100;
        rom[9'b011111_011] = 8'b01000100;
        rom[9'b011111_010] = 8'b01000100;
        rom[9'b011111_001] = 8'b00000000;
        rom[9'b011111_000] = 8'b00000000;

        rom[9'b100000_111] = 8'b00010001;
        rom[9'b100000_110] = 8'b00100010;
        rom[9'b100000_101] = 8'b01000100;
        rom[9'b100000_100] = 8'b10001000;
        rom[9'b100000_011] = 8'b00010001;
        rom[9'b100000_010] = 8'b00100010;
        rom[9'b100000_001] = 8'b01000100;
        rom[9'b100000_000] = 8'b10001000;

        (* font_end *);
    end

endmodule : bitmap_rom
